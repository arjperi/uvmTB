interface top_intf;

    logic [31:0] intf_a;
    logic [31:0] intf_b;
    logic [31:0] intf_c;
    logic intf_clk;
    logic intf_start;

endinterface : top_intf
